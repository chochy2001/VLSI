Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY pwm IS
	--GENERIC(DUTY: INTEGER := 5); -- Ciclo de trabajo
	PORT(DUTY: IN INTEGER RANGE 0 TO 100;
		  CLK1: IN STD_LOGIC;
	     PWM1: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF pwm IS
SIGNAL Q: STD_LOGIC;
SIGNAL CUENTA: INTEGER RANGE 0 TO 100;
BEGIN

	
	PROCESS(CLK1) -- Periodo PWM T = CUENTA/f_CLK
	BEGIN
		IF RISING_EDGE (CLK1) THEN
			IF CUENTA = 100 THEN 
				CUENTA <= 0;
			ELSE 
				CUENTA <= CUENTA + 1;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CUENTA) -- Comparador 
	BEGIN 
		IF CUENTA < DUTY THEN
			Q <= '1';
		ELSE 
			Q <= '0';
		END IF;
	END PROCESS;
		
	PROCESS(CLK1) -- Registro
	BEGIN 
		IF RISING_EDGE(CLK1) THEN
			PWM1 <= Q;
		END IF;
	END PROCESS;
	
END BEAS;