LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY divf IS
	GENERIC(FREC: INTEGER := 249999 ); 
	-- 249999   >> 100 Hz
	-- 24999999 >> 1 Hz
	PORT(CLK_d: IN STD_LOGIC; 
			   CLK: BUFFER STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF divf IS
SIGNAL AUX: INTEGER RANGE 0 TO FREC;
BEGIN
	PROCESS(CLK_d)
	BEGIN
		IF RISING_EDGE (CLK_d) THEN
			IF AUX = 0 THEN
				CLK <= NOT CLK;
				AUX <= FREC;
			ELSE
				AUX <= AUX - 1;
			END IF;
		END IF;
	END PROCESS;

END BEAS;