LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DIVF IS
	GENERIC(FREC: INTEGER := 49999999); -- FREC = (50 MHz/2*Fdeseada) - 1
	-- 24999    >> 1 kHz
	-- 249999   >> 100 Hz
	-- 24999999 >> 1 Hz
	PORT(CLK_MST: IN STD_LOGIC; -- RELOJ PRINCIPAL
			   CLK2: BUFFER STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF DIVF IS
SIGNAL AUX: INTEGER RANGE 0 TO FREC;
BEGIN

	PROCESS(CLK_MST)
	BEGIN
		IF RISING_EDGE (CLK_MST) THEN
			IF AUX = 0 THEN
				CLK2 <= NOT CLK2;
				AUX <= FREC;
			ELSE
				AUX <= AUX - 1;
			END IF;
		END IF;
	END PROCESS;

END BEAS;
