LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DAC IS 
	GENERIC(NBIT: INTEGER:= 7); -- NÚMERO DE BITS DE MI DAC (n-1)
	PORT(CLK, RES: IN STD_LOGIC;
	        DAC_I: IN STD_LOGIC_VECTOR(NBIT DOWNTO 0);
			  DAC_O: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF DAC IS 
SIGNAL DAC_OUT: STD_LOGIC;
SIGNAL DELTA_ADD, SIGMA_ADD, SIGMA_LATCH, DELTA_B: UNSIGNED (NBIT+2 DOWNTO 0);

BEGIN
	DELTA_B (NBIT + 2 DOWNTO NBIT + 1) <= SIGMA_LATCH (NBIT + 2) & SIGMA_LATCH(NBIT + 2);
	DELTA_B (NBIT DOWNTO 0) <= (OTHERS => '0');
	DELTA_ADD <= UNSIGNED ('0' & '0' & DAC_I) + DELTA_B;
	SIGMA_ADD <= DELTA_ADD + SIGMA_LATCH;
	
	PROCESS(CLK, RES)
	BEGIN
		IF RES = '0' THEN
			SIGMA_LATCH <= TO_UNSIGNED (2**(NBIT + 1), SIGMA_LATCH'LENGTH);
			DAC_OUT <= '0';
		ELSIF FALLING_EDGE (CLK) THEN
			SIGMA_LATCH <= SIGMA_ADD;
			DAC_OUT <= SIGMA_LATCH (NBIT + 2);
		END IF;
	END PROCESS;
	
	DAC_O <= DAC_OUT;

END BEAS;