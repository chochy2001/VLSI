LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY Cont IS
	PORT(	CLK: IN STD_LOGIC;
			CUENTA: BUFFER INTEGER RANGE 0 TO 999);
END ENTITY;

ARCHITECTURE BHV of Cont IS
BEGIN
	PROCESS(CLK)
	BEGIN
		IF FALLING_EDGE(CLK) THEN
			IF CUENTA = 999 THEN
				CUENTA <= 0;
			ELSE
				CUENTA <= CUENTA + 1;
			END IF;
		END IF;
	END PROCESS;
END BHV;
			