LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DIVF2 IS
	GENERIC(FREC: INTEGER := 49999999); -- FREC = (50 MHz/2*Fdeseada) - 1
	-- 24999    >> 1 kHz
	-- 249999   >> 100 Hz
	-- 24999999 >> 1 Hz
	PORT(CLK_MST: IN STD_LOGIC; -- RELOJ PRINCIPAL
			   CLK1: BUFFER STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF DIVF2 IS
SIGNAL AUX: INTEGER RANGE 0 TO FREC;
BEGIN

	PROCESS(CLK_MST)
	BEGIN
		IF RISING_EDGE (CLK_MST) THEN
			IF AUX = 0 THEN
				CLK1 <= NOT CLK1;
				AUX <= FREC;
			ELSE
				AUX <= AUX - 1;
			END IF;
		END IF;
	END PROCESS;

END BEAS;